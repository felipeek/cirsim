* Testcase 1
Ve1 1 0 SIN (0 1 0.01meg 0)
Ce8 0 1 3 IC=3m
V1 no3 no2 PWL  (0 1 200u 0.5 500u 2 750u 1 1m 5)
.OP
.TRAN 1u 1m