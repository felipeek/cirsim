* Testcase 1
Ve1 1 0 40
Re2 1 2 10
Ie3 3 2 5
Re4 3 0 10
Re5 2 4 5
Re6 4 0 10
Ge7 0 4 2 4 2
Ce8 0 1 3 IC=3n

.OP
.TRAN 1m 100m