* Testcase 1
* Ve1 1 0 SIN (0 1 0.1meg 0)
* Re2 1 0 3m
Ve1 1 0 SIN(0 9 796 0)
Re2 1 2 30
Le3 2 3 20m
Ce4 3 0 2u
.TRAN 0.00001 0.001