* Testcase 1
Ve1 1 0 SIN (         1   2 3 4          )
Ce8 0 1 3 IC=3m
V1 no3 no2 PWL  (  0 0 5u 3 10u 3 15u 6 40u 6 45u 2 60u 2 65u 0 )
.OP
.TRAN 1m 100m