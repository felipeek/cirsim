* Testcase 1
* Ve1 1 0 SIN (0 1 0.1meg 0)
* Re2 1 0 3m
Ve1 1 0 5
Re2 1 2 1.5
Le3 2 3 10e-3
Ce4 3 0 10e-5
.TRAN 1e-4 1